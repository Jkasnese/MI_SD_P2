`ifndef CHARS
`define CHARS

`define ZERO 8'h30
`define ONE 8'h31
`define TWO  8'h32
`define THREE 8'h33
`define FOUR  8'h34
`define FIVE   8'h35
`define SIX  8'h36
`define SEVEN  8'h37
`define EIGHT  8'h38
`define NINE  8'h39
`define A  8'h41
`define B  8'h42
`define C  8'h43
`define D  8'h44
`define E  8'h45
`define F  8'h46

`endif //CHARS